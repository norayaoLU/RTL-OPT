module mux_dead_mini(
    input x,
    input sel,
    input [7:0] a,        // 8-bit input operand A
    input [7:0] b,        // 8-bit input operand B
    output reg [7:0] result  // Output result
);

// Inline the bitwise operations and combine the logic
always @(*) begin
    if (x) begin
        // And bitwise operation directly
        result = a & b;
    end else begin
        // Or bitwise operation directly
        result = a | b;
    end
end

endmodule