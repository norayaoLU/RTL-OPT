module comparator_8bit (
    input [7:0] A, B,
    output eq, gt, lt
);
    assign eq = (A[7] == B[7]) && (A[6] == B[6]) && (A[5] == B[5]) && (A[4] == B[4]) &&
                (A[3] == B[3]) && (A[2] == B[2]) && (A[1] == B[1]) && (A[0] == B[0]);
    assign gt = (A[7] > B[7]) ||
                ((A[7] == B[7]) && (A[6] > B[6])) ||
                ((A[7] == B[7]) && (A[6] == B[6]) && (A[5] > B[5])) ||
                ((A[7] == B[7]) && (A[6] == B[6]) && (A[5] == B[5]) && (A[4] > B[4])) ||
                ((A[7] == B[7]) && (A[6] == B[6]) && (A[5] == B[5]) && (A[4] == B[4]) && (A[3] > B[3])) ||
                ((A[7] == B[7]) && (A[6] == B[6]) && (A[5] == B[5]) && (A[4] == B[4]) && (A[3] == B[3]) && (A[2] > B[2])) ||
                ((A[7] == B[7]) && (A[6] == B[6]) && (A[5] == B[5]) && (A[4] == B[4]) && (A[3] == B[3]) && (A[2] == B[2]) && (A[1] > B[1])) ||
                ((A[7] == B[7]) && (A[6] == B[6]) && (A[5] == B[5]) && (A[4] == B[4]) && (A[3] == B[3]) && (A[2] == B[2]) && (A[1] == B[1]) && (A[0] > B[0]));
    assign lt = (A[7] < B[7]) ||
                ((A[7] == B[7]) && (A[6] < B[6])) ||
                ((A[7] == B[7]) && (A[6] == B[6]) && (A[5] < B[5])) ||
                ((A[7] == B[7]) && (A[6] == B[6]) && (A[5] == B[5]) && (A[4] < B[4])) ||
                ((A[7] == B[7]) && (A[6] == B[6]) && (A[5] == B[5]) && (A[4] == B[4]) && (A[3] < B[3])) ||
                ((A[7] == B[7]) && (A[6] == B[6]) && (A[5] == B[5]) && (A[4] == B[4]) && (A[3] == B[3]) && (A[2] < B[2])) ||
                ((A[7] == B[7]) && (A[6] == B[6]) && (A[5] == B[5]) && (A[4] == B[4]) && (A[3] == B[3]) && (A[2] == B[2]) && (A[1] < B[1])) ||
                ((A[7] == B[7]) && (A[6] == B[6]) && (A[5] == B[5]) && (A[4] == B[4]) && (A[3] == B[3]) && (A[2] == B[2]) && (A[1] == B[1]) && (A[0] < B[0]));
endmodule