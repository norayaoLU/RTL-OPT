module comparator_4bit (
    input [3:0] A, B,
    output eq, gt, lt
);
    assign eq = (A[3] == B[3]) && (A[2] == B[2]) && (A[1] == B[1]) && (A[0] == B[0]);
    assign gt = (A[3] > B[3]) || 
                ((A[3] == B[3]) && (A[2] > B[2])) || 
                ((A[3] == B[3]) && (A[2] == B[2]) && (A[1] > B[1])) || 
                ((A[3] == B[3]) && (A[2] == B[2]) && (A[1] == B[1]) && (A[0] > B[0]));
    assign lt = (A[3] < B[3]) || 
                ((A[3] == B[3]) && (A[2] < B[2])) || 
                ((A[3] == B[3]) && (A[2] == B[2]) && (A[1] < B[1])) || 
                ((A[3] == B[3]) && (A[2] == B[2]) && (A[1] == B[1]) && (A[0] < B[0]));
endmodule